library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity breakout_game is
	port(
		clk, reset: in std_logic;
		left_btn: in std_logic;
		right_btn: in std_logic;
		vsync: out std_logic;
		hsync: out std_logic;
		state_led: out std_logic_vector(2 downto 0);
		rgb: out std_logic_vector(7 downto 0)
		);
end breakout_game;

architecture arch of breakout_game is
	signal pixel_tick: std_logic;
	signal video_on: std_logic;
	signal pixel_x: std_logic_vector(9 downto 0);
	signal pixel_y: std_logic_vector(9 downto 0);
	
	signal rgb_reg, rgb_next: std_logic_vector(7 downto 0);
	
	signal not_reset, not_left_btn, not_right_btn: std_logic;
	
	type state_type is (newgame, play, newlevel, relevel, over);
	signal state_reg, state_next: state_type;
	
	-- signals used by the number of balls counter
	signal num_balls: std_logic_vector(3 downto 0);
	signal zero_balls: std_logic;
	signal dec_num_balls: std_logic;
	signal clear_num_balls: std_logic;
	
	-- signals used by the level counter
	signal num_levels: std_logic_vector(3 downto 0);
	signal inc_level: std_logic;
	signal clear_level: std_logic;
	
	-- internal status signals generated by the pixel generation circuit
	signal zero_bricks_tick: std_logic;
	signal miss_tick: std_logic;
	
	-- control signals generated by the finite state machine
	signal graph_still: std_logic;
	signal reset_bricks: std_logic;
	
	-- signals used by the timer
	signal timer_tick: std_logic;
	signal timer_done: std_logic;
	signal timer_clear: std_logic;
	
	signal text_on: std_logic_vector(4 downto 0);
	signal graph_on: std_logic_vector(2 downto 0);
	
	signal text_rgb: std_logic_vector(7 downto 0);
	signal graph_rgb: std_logic_vector(7 downto 0);
begin
	-- instantiate the VGA synchronization module
	VGA_sync: entity work.VGA_sync(arch) port map(clk => clk, reset => not_reset,
	video_on => video_on, p_tick => pixel_tick, pixel_x => pixel_x, pixel_y => pixel_y,
	hsync => hsync, vsync => vsync);
	
	-- instantiate the pixel generation module
	pix_gen: entity work.pix_gen_circuit_breakout(arch) port map(clk => clk, reset => not_reset,
	btn => not_left_btn & not_right_btn, video_on => video_on, graph_rgb => graph_rgb, graph_on => graph_on, 
	zero_bricks_tick => zero_bricks_tick, graph_still => graph_still, pixel_x => pixel_x, pixel_y => pixel_y,
	reset_bricks => reset_bricks, miss_tick => miss_tick);

	-- instantiate the text generation module
	text_gen: entity work.text_gen_circuit_breakout(arch) port map(clk => clk, 
	pixel_x => pixel_x, pixel_y => pixel_y, level => num_levels, balls => num_balls, 
	text_on => text_on, text_rgb => text_rgb);
	
	-- instantiate the counter module to count down the number of balls
	ball_counter_unit: entity work.counter(arch) generic map(MIN => 0, MAX => 3, N => 4)
	port map(clk => clk, reset => not_reset, up_down => '1', count => num_balls,
	clear => clear_num_balls, inc_dec => dec_num_balls, zero_flag => zero_balls, full_flag => open);
	
	-- instantiate the counter module to count up the number of levels
	level_counter_unit: entity work.counter(arch) generic map(MIN => 1, MAX => 9, N => 4)
	port map(clk => clk, reset => not_reset, up_down => '0', count => num_levels,
	clear => clear_level, inc_dec => inc_level, zero_flag => open, full_flag => open);
	
	-- instantiate the counter module to implement a timer for the game over screen
	-- the timer_tick signal is asserted at a rate of 60 Hz
	timer_tick <= '1' when pixel_x = "0000000000" and pixel_y = "0000000000" else '0';
	-- to get an 8 second delay implement a counter with an initial value of 480
	timer_unit: entity work.counter(arch) generic map(MIN => 0, MAX => 480, N => 9)
	port map(clk => clk, reset => not_reset, up_down => '1', count => open,
	clear => timer_clear, inc_dec => timer_tick, zero_flag => timer_done, full_flag => open);

	-- take the inverse of the button signals because the push buttons on the Mimas v2 ...
	-- are active low
	not_reset <= not reset;
	not_left_btn <= not left_btn;
	not_right_btn <= not right_btn;
	
	-- registers
	process(clk, not_reset, pixel_tick)
	begin
		if (not_reset = '1') then
			rgb_reg <= (others=>'0');
			state_reg <= newgame;
		elsif (clk'event and clk = '1') then
			if (pixel_tick = '1') then
				rgb_reg <= rgb_next;
			end if;
			state_reg <= state_next;
		end if;
	end process;
	
	-- finite state machine
	process(state_reg, zero_balls, not_left_btn, not_right_btn, miss_tick,
	zero_bricks_tick, timer_done)
	begin
		-- default values
		state_next <= state_reg;
		graph_still <= '1';
		reset_bricks <= '0';
		clear_level <= '0';
		clear_num_balls <= '0';
		inc_level <= '0';
		dec_num_balls <= '0';
		timer_clear <= '0';
		state_led <= "000";
		case state_reg is
			-- in the new game state ...
			when newgame =>
				clear_level <= '1';			-- clear the levels counter
				clear_num_balls <= '1';		-- clear the number of balls counter
				reset_bricks <= '1';			-- reset the bricks
				-- if the player presses any button ...
				if (not_left_btn = '1' or not_right_btn = '1') then
					-- transition into the play state
					state_next <= play;
				end if;
				state_led <= "001";
			-- in the play state ...
			when play =>
				graph_still <= '0';			-- start the animation
				-- if there are no balls left and the player misses the ball ...
				if (zero_balls = '1' and miss_tick = '1') then
					-- transition into the game over state
					state_next <= over;
					timer_clear <= '1';		-- start the count down timer
				-- if the player misses the ball ...
				elsif (miss_tick = '1') then
					dec_num_balls <= '1';	-- decrement the number of balls
					-- transition into the restart level state
					state_next <= relevel;	
				-- if the player clears all the bricks ...
				elsif (zero_bricks_tick = '1') then
					inc_level <= '1';			-- increment the number of levels
					-- transition into the new level state
					state_next <= newlevel;
				end if;
				state_led <= "010";
			-- in the new level state
			when newlevel =>
				reset_bricks <= '1';			-- reset the number of bricks
				-- if the player presses any button ...
				if (not_left_btn = '1' or not_right_btn = '1') then
					-- transition into the play state
					state_next <= play;
				end if;
				state_led <= "011";
			-- in the restart level state
			when relevel =>
				-- if the player presses any button ...
				if (not_left_btn = '1' or not_right_btn = '1') then
					-- transition into the play state
					state_next <= play;
				end if;
				state_led <= "100";
			-- in the game over state
			when over =>
				-- wait until the timer is finished ...
				if (timer_done = '1') then
					-- then transition into the new game state
					state_next <= newgame;
				end if;
				state_led <= "101";
		end case;
	end process;
	
	-- rgb multiplexing circuit
	process(video_on, graph_on, text_on, text_rgb, graph_rgb, state_reg)
	begin
		-- if in the border area of the screen ...
		if (video_on = '0') then
			-- set the pixel color to black
			rgb_next <= (others=>'0');
		-- if in the display area of the screen ...
		else
			-- display the game objects
			-- the priority in the if-else statement determines whether the object is in the foreground or the background
			-- if in the new game or game over states ...
			if (state_reg = newgame and (text_on(1) = '1' or text_on(2) = '1')) or
				(state_reg = over and (text_on(0) = '1')) then
				-- give priority to the text objects so the name, game over message and rules are in the foreground
				rgb_next <= text_rgb;
			elsif (graph_on /= "000") then
				rgb_next <= graph_rgb;
			elsif (text_on(3) = '1' or text_on(4) = '1') then
				rgb_next <= text_rgb;
			else
				-- background color
				rgb_next <= "11111100";
			end if;
		end if;
	end process;
	
	rgb <= rgb_reg;
	
end arch;

